interface intf();
   logic a;
   logic b;
   logic c;
   logic sum;
   logic carry;
  
endinterface
