----------------Generation of values-----------
# a=1 b=1 c=0 sum=0 carry=0
# ----------------Generation of values-----------
# a=0 b=1 c=1 sum=0 carry=0
# ----------------Generation of values-----------
# a=1 b=1 c=0 sum=0 carry=0
# ----------------received values of trans-----------
# a=0 b=0 c=1 sum=0 carry=0
# ----------------monitor received-----------
# a=0 b=0 c=1 sum=1 carry=0
# ----------------scoreboard received-----------
# a=0 b=0 c=1 sum=1 carry=0
# -----------------pass-------------
# -------------transaction done--------
# 
# ----------------received values of trans-----------
# a=0 b=0 c=1 sum=0 carry=0
# ----------------monitor received-----------
# a=0 b=0 c=1 sum=1 carry=0
# ----------------scoreboard received-----------
# a=0 b=0 c=1 sum=1 carry=0
# -----------------pass-------------
# -------------transaction done--------
# 
# ----------------received values of trans-----------
# a=0 b=0 c=1 sum=0 carry=0
# ----------------monitor received-----------
# a=0 b=0 c=1 sum=1 carry=0
# ----------------scoreboard received-----------
# a=0 b=0 c=1 sum=1 carry=0
# -----------------pass-------------
# -------------transaction done--------
